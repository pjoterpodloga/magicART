magic
tech scmos
timestamp 1700319599
<< nwell >>
rect 23 141 252 222
<< electrodecontact >>
rect 197 107 202 112
rect 197 97 202 102
rect 197 87 202 92
rect 197 77 202 82
<< electrodecap >>
rect 194 67 243 118
rect 154 14 243 67
<< ntransistor >>
rect 51 93 56 118
rect 67 93 72 118
rect 83 93 88 118
rect 99 93 104 118
rect 115 93 120 118
rect 131 93 136 118
rect 147 93 152 118
rect 163 93 168 118
rect 51 44 56 62
rect 67 44 72 62
rect 83 44 88 62
rect 99 44 104 62
rect 115 44 120 62
rect 131 44 136 62
rect 51 15 56 33
rect 67 15 72 33
rect 83 15 88 33
rect 99 15 104 33
rect 115 15 120 33
rect 131 15 136 33
<< ptransistor >>
rect 43 189 48 207
rect 83 189 88 207
rect 99 189 104 207
rect 115 189 120 207
rect 131 189 136 207
rect 147 189 152 207
rect 163 189 168 207
rect 179 189 184 207
rect 195 189 200 207
rect 211 189 216 207
rect 227 189 232 207
rect 43 160 48 178
rect 83 160 88 178
rect 99 160 104 178
rect 115 160 120 178
rect 131 160 136 178
rect 147 160 152 178
rect 163 160 168 178
rect 179 160 184 178
rect 195 160 200 178
rect 211 160 216 178
rect 227 160 232 178
rect 43 147 48 152
<< ndiffusion >>
rect 48 93 51 118
rect 56 93 59 118
rect 64 93 67 118
rect 72 93 75 118
rect 80 93 83 118
rect 88 93 91 118
rect 96 93 99 118
rect 104 93 107 118
rect 112 93 115 118
rect 120 93 123 118
rect 128 93 131 118
rect 136 93 139 118
rect 144 93 147 118
rect 152 93 155 118
rect 160 93 163 118
rect 168 93 171 118
rect 48 44 51 62
rect 56 44 59 62
rect 64 44 67 62
rect 72 44 75 62
rect 80 44 83 62
rect 88 44 91 62
rect 96 44 99 62
rect 104 44 107 62
rect 112 44 115 62
rect 120 44 123 62
rect 128 44 131 62
rect 136 44 139 62
rect 48 15 51 33
rect 56 15 59 33
rect 64 15 67 33
rect 72 15 75 33
rect 80 15 83 33
rect 88 15 91 33
rect 96 15 99 33
rect 104 15 107 33
rect 112 15 115 33
rect 120 15 123 33
rect 128 15 131 33
rect 136 15 139 33
<< pdiffusion >>
rect 40 189 43 207
rect 48 189 51 207
rect 80 189 83 207
rect 88 189 91 207
rect 96 189 99 207
rect 104 189 107 207
rect 112 189 115 207
rect 120 189 123 207
rect 128 189 131 207
rect 136 189 139 207
rect 144 189 147 207
rect 152 189 155 207
rect 160 189 163 207
rect 168 189 171 207
rect 176 189 179 207
rect 184 189 187 207
rect 192 189 195 207
rect 200 189 203 207
rect 208 189 211 207
rect 216 189 219 207
rect 224 189 227 207
rect 232 189 235 207
rect 40 160 43 178
rect 48 160 51 178
rect 80 160 83 178
rect 88 160 91 178
rect 96 160 99 178
rect 104 160 107 178
rect 112 160 115 178
rect 120 160 123 178
rect 128 160 131 178
rect 136 160 139 178
rect 144 160 147 178
rect 152 160 155 178
rect 160 160 163 178
rect 168 160 171 178
rect 176 160 179 178
rect 184 160 187 178
rect 192 160 195 178
rect 200 160 203 178
rect 208 160 211 178
rect 216 160 219 178
rect 224 160 227 178
rect 232 160 235 178
rect 40 147 43 152
rect 48 147 51 152
<< ndcontact >>
rect 43 93 48 118
rect 59 93 64 118
rect 75 93 80 118
rect 91 93 96 118
rect 107 93 112 118
rect 123 93 128 118
rect 139 93 144 118
rect 155 93 160 118
rect 171 93 176 118
rect 43 44 48 62
rect 59 44 64 62
rect 75 44 80 62
rect 91 44 96 62
rect 107 44 112 62
rect 123 44 128 62
rect 139 44 144 62
rect 43 15 48 33
rect 59 15 64 33
rect 75 15 80 33
rect 91 15 96 33
rect 107 15 112 33
rect 123 15 128 33
rect 139 15 144 33
<< pdcontact >>
rect 35 189 40 207
rect 51 189 56 207
rect 75 189 80 207
rect 91 189 96 207
rect 107 189 112 207
rect 123 189 128 207
rect 139 189 144 207
rect 155 189 160 207
rect 171 189 176 207
rect 187 189 192 207
rect 203 189 208 207
rect 219 189 224 207
rect 235 189 240 207
rect 35 160 40 178
rect 51 160 56 178
rect 75 160 80 178
rect 91 160 96 178
rect 107 160 112 178
rect 123 160 128 178
rect 139 160 144 178
rect 155 160 160 178
rect 171 160 176 178
rect 187 160 192 178
rect 203 160 208 178
rect 219 160 224 178
rect 235 160 240 178
rect 35 147 40 152
rect 51 147 56 152
<< psubstratepcontact >>
rect 11 229 16 234
rect 27 229 32 234
rect 43 229 48 234
rect 59 229 64 234
rect 75 229 80 234
rect 91 229 96 234
rect 107 229 112 234
rect 123 229 128 234
rect 139 229 144 234
rect 155 229 160 234
rect 171 229 176 234
rect 187 229 192 234
rect 203 229 208 234
rect 219 229 224 234
rect 235 229 240 234
rect 251 229 256 234
rect 1 219 6 224
rect 260 219 265 224
rect 1 203 6 208
rect 1 187 6 192
rect 260 203 265 208
rect 260 187 265 192
rect 1 171 6 176
rect 1 155 6 160
rect 260 171 265 176
rect 260 155 265 160
rect 1 139 6 144
rect 260 139 265 144
rect 1 123 6 128
rect 260 123 265 128
rect 1 107 6 112
rect 1 91 6 96
rect 260 107 265 112
rect 260 91 265 96
rect 1 75 6 80
rect 260 75 265 80
rect 1 59 6 64
rect 1 43 6 48
rect 1 27 6 32
rect 1 11 6 16
rect 260 59 265 64
rect 260 43 265 48
rect 260 27 265 32
rect 260 11 265 16
rect 11 1 16 6
rect 27 1 32 6
rect 43 1 48 6
rect 59 1 64 6
rect 75 1 80 6
rect 91 1 96 6
rect 107 1 112 6
rect 123 1 128 6
rect 139 1 144 6
rect 155 1 160 6
rect 171 1 176 6
rect 187 1 192 6
rect 203 1 208 6
rect 219 1 224 6
rect 235 1 240 6
rect 250 1 255 6
<< nsubstratencontact >>
rect 35 214 40 219
rect 45 214 50 219
rect 55 214 60 219
rect 65 214 70 219
rect 75 214 80 219
rect 86 214 91 219
rect 96 214 101 219
rect 107 214 112 219
rect 118 214 123 219
rect 128 214 133 219
rect 139 214 144 219
rect 150 214 155 219
rect 160 214 165 219
rect 171 214 176 219
rect 182 214 187 219
rect 192 214 197 219
rect 203 214 208 219
rect 214 214 219 219
rect 224 214 229 219
rect 235 214 240 219
rect 26 208 31 213
rect 26 198 31 203
rect 26 188 31 193
rect 244 205 249 210
rect 244 194 249 199
rect 26 178 31 183
rect 244 183 249 188
rect 26 168 31 173
rect 26 158 31 163
rect 244 172 249 177
rect 244 161 249 166
rect 26 148 31 153
rect 244 150 249 155
<< polysilicon >>
rect 43 207 48 210
rect 83 207 88 210
rect 99 207 104 210
rect 115 207 120 210
rect 131 207 136 210
rect 147 207 152 210
rect 163 207 168 210
rect 179 207 184 210
rect 195 207 200 210
rect 211 207 216 210
rect 227 207 232 210
rect 43 186 48 189
rect 83 186 88 189
rect 99 186 104 189
rect 115 186 120 189
rect 131 186 136 189
rect 147 186 152 189
rect 163 186 168 189
rect 179 186 184 189
rect 195 186 200 189
rect 211 186 216 189
rect 227 186 232 189
rect 43 181 51 186
rect 83 181 232 186
rect 43 178 48 181
rect 83 178 88 181
rect 99 178 104 181
rect 115 178 120 181
rect 131 178 136 181
rect 147 178 152 181
rect 163 178 168 181
rect 179 178 184 181
rect 195 178 200 181
rect 211 178 216 181
rect 227 178 232 181
rect 43 158 48 160
rect 83 157 88 160
rect 99 157 104 160
rect 115 157 120 160
rect 131 157 136 160
rect 43 152 48 154
rect 147 147 152 160
rect 163 157 168 160
rect 179 157 184 160
rect 195 157 200 160
rect 211 157 216 160
rect 227 157 232 160
rect 43 142 48 147
rect 30 123 168 128
rect 51 118 56 123
rect 67 118 72 120
rect 83 118 88 120
rect 99 118 104 123
rect 115 118 120 123
rect 131 118 136 120
rect 147 118 152 120
rect 163 118 168 123
rect 182 112 248 123
rect 182 107 184 112
rect 189 107 248 112
rect 182 102 248 107
rect 182 97 184 102
rect 189 97 248 102
rect 51 91 56 93
rect 67 88 72 93
rect 83 88 88 93
rect 99 91 104 93
rect 115 91 120 93
rect 131 88 136 93
rect 147 88 152 93
rect 163 91 168 93
rect 182 92 248 97
rect 30 83 152 88
rect 182 87 184 92
rect 189 87 248 92
rect 182 72 248 87
rect 51 62 56 64
rect 67 62 72 64
rect 83 62 88 64
rect 99 62 104 64
rect 115 62 120 64
rect 131 62 136 64
rect 51 41 56 44
rect 67 41 72 44
rect 83 41 88 44
rect 99 41 104 44
rect 115 41 120 44
rect 131 41 136 44
rect 48 36 136 41
rect 51 33 56 36
rect 67 33 72 36
rect 83 33 88 36
rect 99 33 104 36
rect 115 33 120 36
rect 131 33 136 36
rect 51 13 56 15
rect 67 13 72 15
rect 83 13 88 15
rect 99 13 104 15
rect 115 13 120 15
rect 131 13 136 15
rect 149 9 248 72
<< polycontact >>
rect 51 181 56 186
rect 147 142 152 147
rect 43 137 48 142
rect 184 107 189 112
rect 184 97 189 102
rect 184 87 189 92
rect 35 36 48 41
<< metal1 >>
rect 0 234 266 235
rect 0 229 11 234
rect 16 229 27 234
rect 32 229 43 234
rect 48 229 59 234
rect 64 229 75 234
rect 80 229 91 234
rect 96 229 107 234
rect 112 229 123 234
rect 128 229 139 234
rect 144 229 155 234
rect 160 229 171 234
rect 176 229 187 234
rect 192 229 203 234
rect 208 229 219 234
rect 224 229 235 234
rect 240 229 251 234
rect 256 229 266 234
rect 0 228 266 229
rect 0 224 7 228
rect 0 219 1 224
rect 6 219 7 224
rect 259 224 266 228
rect 0 208 7 219
rect 0 203 1 208
rect 6 203 7 208
rect 0 192 7 203
rect 0 187 1 192
rect 6 187 7 192
rect 0 176 7 187
rect 0 171 1 176
rect 6 171 7 176
rect 0 160 7 171
rect 0 155 1 160
rect 6 155 7 160
rect 0 144 7 155
rect 25 219 250 220
rect 25 214 35 219
rect 40 214 45 219
rect 50 214 55 219
rect 60 214 65 219
rect 70 214 75 219
rect 80 214 86 219
rect 91 214 96 219
rect 101 214 107 219
rect 112 214 118 219
rect 123 214 128 219
rect 133 214 139 219
rect 144 214 150 219
rect 155 214 160 219
rect 165 214 171 219
rect 176 214 182 219
rect 187 214 192 219
rect 197 214 203 219
rect 208 214 214 219
rect 219 214 224 219
rect 229 214 235 219
rect 240 214 250 219
rect 25 213 250 214
rect 25 208 26 213
rect 31 208 32 213
rect 25 203 32 208
rect 25 198 26 203
rect 31 198 32 203
rect 25 193 32 198
rect 25 188 26 193
rect 31 188 32 193
rect 25 183 32 188
rect 25 178 26 183
rect 31 178 32 183
rect 25 173 32 178
rect 25 168 26 173
rect 31 168 32 173
rect 25 163 32 168
rect 25 158 26 163
rect 31 158 32 163
rect 25 153 32 158
rect 25 148 26 153
rect 31 148 32 153
rect 25 147 32 148
rect 35 207 40 213
rect 75 207 80 213
rect 107 207 112 213
rect 139 207 144 213
rect 171 207 176 213
rect 203 207 208 213
rect 235 207 240 213
rect 56 189 72 207
rect 35 178 40 189
rect 51 178 56 181
rect 56 160 64 178
rect 35 152 40 160
rect 0 139 1 144
rect 6 139 7 144
rect 51 142 56 147
rect 0 128 7 139
rect 0 123 1 128
rect 6 123 7 128
rect 0 112 7 123
rect 0 107 1 112
rect 6 107 7 112
rect 0 96 7 107
rect 0 91 1 96
rect 6 91 7 96
rect 0 80 7 91
rect 0 75 1 80
rect 6 75 7 80
rect 0 64 7 75
rect 0 59 1 64
rect 6 59 7 64
rect 0 48 7 59
rect 0 43 1 48
rect 6 43 7 48
rect 0 32 7 43
rect 35 137 43 142
rect 48 137 56 142
rect 35 41 40 137
rect 59 134 64 160
rect 67 147 72 189
rect 75 178 80 189
rect 91 178 96 189
rect 107 178 112 189
rect 123 178 128 189
rect 139 178 144 189
rect 155 178 160 189
rect 171 178 176 189
rect 187 178 192 189
rect 203 178 208 189
rect 219 178 224 189
rect 235 178 240 189
rect 243 210 250 213
rect 243 205 244 210
rect 249 205 250 210
rect 243 199 250 205
rect 243 194 244 199
rect 249 194 250 199
rect 243 188 250 194
rect 243 183 244 188
rect 249 183 250 188
rect 243 177 250 183
rect 243 172 244 177
rect 249 172 250 177
rect 243 166 250 172
rect 243 161 244 166
rect 249 161 250 166
rect 91 157 96 160
rect 123 157 128 160
rect 155 157 160 160
rect 187 157 192 160
rect 219 157 224 160
rect 91 152 224 157
rect 243 155 250 161
rect 67 142 147 147
rect 152 142 189 147
rect 43 129 176 134
rect 43 118 48 129
rect 59 121 96 126
rect 59 118 64 121
rect 91 118 96 121
rect 59 70 64 93
rect 75 82 80 93
rect 107 118 112 129
rect 123 121 160 126
rect 123 118 128 121
rect 155 118 160 121
rect 91 90 96 93
rect 123 90 128 93
rect 91 85 128 90
rect 171 118 176 129
rect 184 112 189 142
rect 184 102 189 107
rect 139 82 144 93
rect 184 92 189 97
rect 184 82 189 87
rect 75 77 189 82
rect 197 126 202 152
rect 243 150 244 155
rect 249 150 250 155
rect 243 149 250 150
rect 259 219 260 224
rect 265 219 266 224
rect 259 208 266 219
rect 259 203 260 208
rect 265 203 266 208
rect 259 192 266 203
rect 259 187 260 192
rect 265 187 266 192
rect 259 176 266 187
rect 259 171 260 176
rect 265 171 266 176
rect 259 160 266 171
rect 259 155 260 160
rect 265 155 266 160
rect 259 144 266 155
rect 259 139 260 144
rect 265 139 266 144
rect 259 128 266 139
rect 197 121 239 126
rect 259 123 260 128
rect 265 123 266 128
rect 197 112 202 121
rect 197 102 202 107
rect 197 92 202 97
rect 197 82 202 87
rect 197 72 202 77
rect 43 65 64 70
rect 75 68 202 72
rect 259 112 266 123
rect 259 107 260 112
rect 265 107 266 112
rect 259 96 266 107
rect 259 91 260 96
rect 265 91 266 96
rect 259 80 266 91
rect 259 75 260 80
rect 265 75 266 80
rect 75 67 144 68
rect 43 62 48 65
rect 75 62 80 67
rect 107 62 112 67
rect 139 62 144 67
rect 0 27 1 32
rect 6 27 7 32
rect 0 16 7 27
rect 0 11 1 16
rect 6 11 7 16
rect 43 33 48 36
rect 59 33 64 44
rect 75 33 80 44
rect 91 33 96 44
rect 107 33 112 44
rect 123 33 128 44
rect 139 33 144 44
rect 259 64 266 75
rect 259 59 260 64
rect 265 59 266 64
rect 259 48 266 59
rect 259 43 260 48
rect 265 43 266 48
rect 259 32 266 43
rect 259 27 260 32
rect 265 27 266 32
rect 259 16 266 27
rect 0 7 7 11
rect 59 7 64 15
rect 91 7 96 15
rect 123 7 128 15
rect 259 11 260 16
rect 265 11 266 16
rect 259 7 266 11
rect 0 6 266 7
rect 0 1 11 6
rect 16 1 27 6
rect 32 1 43 6
rect 48 1 59 6
rect 64 1 75 6
rect 80 1 91 6
rect 96 1 107 6
rect 112 1 123 6
rect 128 1 139 6
rect 144 1 155 6
rect 160 1 171 6
rect 176 1 187 6
rect 192 1 203 6
rect 208 1 219 6
rect 224 1 235 6
rect 240 1 250 6
rect 255 1 266 6
rect 0 0 266 1
<< labels >>
rlabel metal1 139 15 144 62 1 out
rlabel metal1 107 15 112 62 1 out
rlabel metal1 75 15 80 62 1 out
rlabel metal1 123 15 128 62 1 Gnd
rlabel metal1 91 15 96 62 1 Gnd
rlabel metal1 59 15 64 62 1 Gnd
rlabel polysilicon 30 123 35 128 4 inn
rlabel polysilicon 30 83 35 88 2 inp
rlabel metal1 234 121 239 126 1 out
rlabel nwell 35 214 240 219 1 Vdd
rlabel ndcontact 43 15 48 33 1 4
rlabel ndcontact 43 44 48 62 1 3
rlabel ndcontact 59 93 64 118 1 3
rlabel ndcontact 91 93 96 118 1 3
rlabel ndcontact 123 93 128 118 1 3
rlabel ndcontact 155 93 160 118 1 3
rlabel ndcontact 171 93 176 118 1 1
rlabel ndcontact 139 93 144 118 1 2
<< end >>
